module control_unit (
    input wire clk,
    input wire reset,

    //Instruction

    //Flags

    //Mux controllers

    //Register controllers
    
    //Functional controllers
);
    
    //State and cycle variables

    //Parameters
        //States
        //Opcodes
        //Other parameters

    //Startup handler

    //Transition function

    //State output handler
endmodule