module cpu_MIPS (
    input wire clk,
    input wire reset
);

// Control wires

// Data wires

// Flag wires

// Instantiating modules

    //Muxes

    //Registers

    //Provided modules

    //Miscellaneous modules

    //Control unit

endmodule