module cpu_MIPS (
    input wire clk,
    input wire reset
);

// Control wires

// Data wires

// Flag wires

// Instantiating modules

endmodule